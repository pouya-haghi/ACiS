`timescale 1ns / 1ps


module runtimeLoadtable(
    input logic clk, 
    input logic rst,
    input logic [dwidth_RFadd-1:0] wr_add,
    input logic [num_col-1:0] wr_en,
    input logic [phit_size-1:0] wr_data
    );
    
    
endmodule
