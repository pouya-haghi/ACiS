`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/10/2021 05:59:24 PM
// Design Name: 
// Module Name: package_mine
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
package package_mine;
//    interface data_channel;
//    logic [63:0] inp1, inp2, out1;
//    endinterface

//    interface control_channel;
//    logic [1:0] op;
//    endinterface
    typedef enum {ADD, SUB} op_list;
endpackage
