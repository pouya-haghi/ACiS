parameter tb_fifo_width=32;
parameter tb_fifo_size=5;