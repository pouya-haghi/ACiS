interface data_channel;
logic [63:0] inp1, inp2, out1;
endinterface

interface control_channel;
logic [1:0] op;
endinterface