`timescale 1ns / 1ps

module float_generator(
    input  logic [4:0] count,
    output logic [31:0] float
    );
    
    always_comb begin
    case(count)
        5'b00000: float = 32'b00000000000000000000000000000000;
        5'b00001: float = 32'b00111111100000000000000000000000;
        5'b00010: float = 32'b01000000000000000000000000000000;
        5'b00011: float = 32'b01000000010000000000000000000000;
        5'b00100: float = 32'b01000000100000000000000000000000;
        5'b00101: float = 32'b01000000101000000000000000000000;
        5'b00110: float = 32'b01000000110000000000000000000000; 
        5'b00111: float = 32'b01000000111000000000000000000000;
        5'b01000: float = 32'b01000001000000000000000000000000;
        5'b01001: float = 32'b01000001000100000000000000000000;
        5'b01010: float = 32'b01000001001000000000000000000000;
        5'b01011: float = 32'b01000001001100000000000000000000;
        5'b01100: float = 32'b01000001010000000000000000000000;
        5'b01101: float = 32'b01000001010100000000000000000000;
        5'b01110: float = 32'b01000001011000000000000000000000;
        5'b01111: float = 32'b01000001011100000000000000000000;
        5'b10000: float = 32'b01000001100000000000000000000000;
        5'b10001: float = 32'b01000001100010000000000000000000;
        5'b10010: float = 32'b01000001100100000000000000000000;
        5'b10011: float = 32'b01000001100110000000000000000000;
        5'b10100: float = 32'b01000001101000000000000000000000;
        5'b10101: float = 32'b01000001101010000000000000000000;
        5'b10110: float = 32'b01000001101100000000000000000000;
        5'b10111: float = 32'b01000001101110000000000000000000;
        5'b11000: float = 32'b01000001110000000000000000000000;
        5'b11001: float = 32'b01000001110010000000000000000000;
        5'b11010: float = 32'b01000001110100000000000000000000;
        5'b11011: float = 32'b01000001110110000000000000000000;
        5'b11100: float = 32'b01000001111000000000000000000000;
        5'b11101: float = 32'b01000001111010000000000000000000;
        5'b11110: float = 32'b01000001111100000000000000000000;
        5'b11111: float = 32'b01000001111110000000000000000000;
        default:  float = 32'b00000000000000000000000000000000;
    endcase
    end
endmodule
